
module top();
   logic [7:0] data;
   logic [15:0] addr;
   logic 	rst_l; 
   logic 	clock_15;
   logic 	sndirq, sndnmi;

   //Block RAM for system memory

   
   //Block ROM for program memory

   
   //6502 Processor Instantiation

   
   //Pokey Audio Synthesis Chip

   
   //PWM Audio output interface

   
   
endmodule: top
